`include "cash.v"

module FastMult(
    input wire[3:0] io_lhs,
    input wire[3:0] io_rhs,
    output wire[7:0] io_out
);
    reg[7:0] m10[0:255];
    wire[7:0] w13, w15, a17, a18;

    initial begin
        m10[0] = 8'h0;
        m10[1] = 8'h0;
        m10[2] = 8'h0;
        m10[3] = 8'h0;
        m10[4] = 8'h0;
        m10[5] = 8'h0;
        m10[6] = 8'h0;
        m10[7] = 8'h0;
        m10[8] = 8'h0;
        m10[9] = 8'h0;
        m10[10] = 8'h0;
        m10[11] = 8'h0;
        m10[12] = 8'h0;
        m10[13] = 8'h0;
        m10[14] = 8'h0;
        m10[15] = 8'h0;
        m10[16] = 8'h0;
        m10[17] = 8'h1;
        m10[18] = 8'h2;
        m10[19] = 8'h3;
        m10[20] = 8'h4;
        m10[21] = 8'h5;
        m10[22] = 8'h6;
        m10[23] = 8'h7;
        m10[24] = 8'h8;
        m10[25] = 8'h9;
        m10[26] = 8'ha;
        m10[27] = 8'hb;
        m10[28] = 8'hc;
        m10[29] = 8'hd;
        m10[30] = 8'he;
        m10[31] = 8'hf;
        m10[32] = 8'h0;
        m10[33] = 8'h2;
        m10[34] = 8'h4;
        m10[35] = 8'h6;
        m10[36] = 8'h8;
        m10[37] = 8'ha;
        m10[38] = 8'hc;
        m10[39] = 8'he;
        m10[40] = 8'h10;
        m10[41] = 8'h12;
        m10[42] = 8'h14;
        m10[43] = 8'h16;
        m10[44] = 8'h18;
        m10[45] = 8'h1a;
        m10[46] = 8'h1c;
        m10[47] = 8'h1e;
        m10[48] = 8'h0;
        m10[49] = 8'h3;
        m10[50] = 8'h6;
        m10[51] = 8'h9;
        m10[52] = 8'hc;
        m10[53] = 8'hf;
        m10[54] = 8'h12;
        m10[55] = 8'h15;
        m10[56] = 8'h18;
        m10[57] = 8'h1b;
        m10[58] = 8'h1e;
        m10[59] = 8'h21;
        m10[60] = 8'h24;
        m10[61] = 8'h27;
        m10[62] = 8'h2a;
        m10[63] = 8'h2d;
        m10[64] = 8'h0;
        m10[65] = 8'h4;
        m10[66] = 8'h8;
        m10[67] = 8'hc;
        m10[68] = 8'h10;
        m10[69] = 8'h14;
        m10[70] = 8'h18;
        m10[71] = 8'h1c;
        m10[72] = 8'h20;
        m10[73] = 8'h24;
        m10[74] = 8'h28;
        m10[75] = 8'h2c;
        m10[76] = 8'h30;
        m10[77] = 8'h34;
        m10[78] = 8'h38;
        m10[79] = 8'h3c;
        m10[80] = 8'h0;
        m10[81] = 8'h5;
        m10[82] = 8'ha;
        m10[83] = 8'hf;
        m10[84] = 8'h14;
        m10[85] = 8'h19;
        m10[86] = 8'h1e;
        m10[87] = 8'h23;
        m10[88] = 8'h28;
        m10[89] = 8'h2d;
        m10[90] = 8'h32;
        m10[91] = 8'h37;
        m10[92] = 8'h3c;
        m10[93] = 8'h41;
        m10[94] = 8'h46;
        m10[95] = 8'h4b;
        m10[96] = 8'h0;
        m10[97] = 8'h6;
        m10[98] = 8'hc;
        m10[99] = 8'h12;
        m10[100] = 8'h18;
        m10[101] = 8'h1e;
        m10[102] = 8'h24;
        m10[103] = 8'h2a;
        m10[104] = 8'h30;
        m10[105] = 8'h36;
        m10[106] = 8'h3c;
        m10[107] = 8'h42;
        m10[108] = 8'h48;
        m10[109] = 8'h4e;
        m10[110] = 8'h54;
        m10[111] = 8'h5a;
        m10[112] = 8'h0;
        m10[113] = 8'h7;
        m10[114] = 8'he;
        m10[115] = 8'h15;
        m10[116] = 8'h1c;
        m10[117] = 8'h23;
        m10[118] = 8'h2a;
        m10[119] = 8'h31;
        m10[120] = 8'h38;
        m10[121] = 8'h3f;
        m10[122] = 8'h46;
        m10[123] = 8'h4d;
        m10[124] = 8'h54;
        m10[125] = 8'h5b;
        m10[126] = 8'h62;
        m10[127] = 8'h69;
        m10[128] = 8'h0;
        m10[129] = 8'h8;
        m10[130] = 8'h10;
        m10[131] = 8'h18;
        m10[132] = 8'h20;
        m10[133] = 8'h28;
        m10[134] = 8'h30;
        m10[135] = 8'h38;
        m10[136] = 8'h40;
        m10[137] = 8'h48;
        m10[138] = 8'h50;
        m10[139] = 8'h58;
        m10[140] = 8'h60;
        m10[141] = 8'h68;
        m10[142] = 8'h70;
        m10[143] = 8'h78;
        m10[144] = 8'h0;
        m10[145] = 8'h9;
        m10[146] = 8'h12;
        m10[147] = 8'h1b;
        m10[148] = 8'h24;
        m10[149] = 8'h2d;
        m10[150] = 8'h36;
        m10[151] = 8'h3f;
        m10[152] = 8'h48;
        m10[153] = 8'h51;
        m10[154] = 8'h5a;
        m10[155] = 8'h63;
        m10[156] = 8'h6c;
        m10[157] = 8'h75;
        m10[158] = 8'h7e;
        m10[159] = 8'h87;
        m10[160] = 8'h0;
        m10[161] = 8'ha;
        m10[162] = 8'h14;
        m10[163] = 8'h1e;
        m10[164] = 8'h28;
        m10[165] = 8'h32;
        m10[166] = 8'h3c;
        m10[167] = 8'h46;
        m10[168] = 8'h50;
        m10[169] = 8'h5a;
        m10[170] = 8'h64;
        m10[171] = 8'h6e;
        m10[172] = 8'h78;
        m10[173] = 8'h82;
        m10[174] = 8'h8c;
        m10[175] = 8'h96;
        m10[176] = 8'h0;
        m10[177] = 8'hb;
        m10[178] = 8'h16;
        m10[179] = 8'h21;
        m10[180] = 8'h2c;
        m10[181] = 8'h37;
        m10[182] = 8'h42;
        m10[183] = 8'h4d;
        m10[184] = 8'h58;
        m10[185] = 8'h63;
        m10[186] = 8'h6e;
        m10[187] = 8'h79;
        m10[188] = 8'h84;
        m10[189] = 8'h8f;
        m10[190] = 8'h9a;
        m10[191] = 8'ha5;
        m10[192] = 8'h0;
        m10[193] = 8'hc;
        m10[194] = 8'h18;
        m10[195] = 8'h24;
        m10[196] = 8'h30;
        m10[197] = 8'h3c;
        m10[198] = 8'h48;
        m10[199] = 8'h54;
        m10[200] = 8'h60;
        m10[201] = 8'h6c;
        m10[202] = 8'h78;
        m10[203] = 8'h84;
        m10[204] = 8'h90;
        m10[205] = 8'h9c;
        m10[206] = 8'ha8;
        m10[207] = 8'hb4;
        m10[208] = 8'h0;
        m10[209] = 8'hd;
        m10[210] = 8'h1a;
        m10[211] = 8'h27;
        m10[212] = 8'h34;
        m10[213] = 8'h41;
        m10[214] = 8'h4e;
        m10[215] = 8'h5b;
        m10[216] = 8'h68;
        m10[217] = 8'h75;
        m10[218] = 8'h82;
        m10[219] = 8'h8f;
        m10[220] = 8'h9c;
        m10[221] = 8'ha9;
        m10[222] = 8'hb6;
        m10[223] = 8'hc3;
        m10[224] = 8'h0;
        m10[225] = 8'he;
        m10[226] = 8'h1c;
        m10[227] = 8'h2a;
        m10[228] = 8'h38;
        m10[229] = 8'h46;
        m10[230] = 8'h54;
        m10[231] = 8'h62;
        m10[232] = 8'h70;
        m10[233] = 8'h7e;
        m10[234] = 8'h8c;
        m10[235] = 8'h9a;
        m10[236] = 8'ha8;
        m10[237] = 8'hb6;
        m10[238] = 8'hc4;
        m10[239] = 8'hd2;
        m10[240] = 8'h0;
        m10[241] = 8'hf;
        m10[242] = 8'h1e;
        m10[243] = 8'h2d;
        m10[244] = 8'h3c;
        m10[245] = 8'h4b;
        m10[246] = 8'h5a;
        m10[247] = 8'h69;
        m10[248] = 8'h78;
        m10[249] = 8'h87;
        m10[250] = 8'h96;
        m10[251] = 8'ha5;
        m10[252] = 8'hb4;
        m10[253] = 8'hc3;
        m10[254] = 8'hd2;
        m10[255] = 8'he1;
    end
    assign w13 = {4'h0, io_rhs};
    assign w15 = {4'h0, io_lhs};
    assign a17 = w15 << 8'h4;
    assign a18 = a17 | w13;

    assign io_out = m10[a18];

endmodule
