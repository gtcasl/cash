module FastMult(
  input wire[3:0] io_lhs,
  input wire[3:0] io_rhs,
  output wire[7:0] io_out
);
  reg[7:0] mem8[0:255]; // fastmult.cpp(20)
  wire[7:0] zext9;
  wire[7:0] zext11;
  wire[7:0] sll15;
  wire[7:0] or17;

  initial begin
    mem8[0] = 8'h0;
    mem8[1] = 8'h0;
    mem8[2] = 8'h0;
    mem8[3] = 8'h0;
    mem8[4] = 8'h0;
    mem8[5] = 8'h0;
    mem8[6] = 8'h0;
    mem8[7] = 8'h0;
    mem8[8] = 8'h0;
    mem8[9] = 8'h0;
    mem8[10] = 8'h0;
    mem8[11] = 8'h0;
    mem8[12] = 8'h0;
    mem8[13] = 8'h0;
    mem8[14] = 8'h0;
    mem8[15] = 8'h0;
    mem8[16] = 8'h0;
    mem8[17] = 8'h1;
    mem8[18] = 8'h2;
    mem8[19] = 8'h3;
    mem8[20] = 8'h4;
    mem8[21] = 8'h5;
    mem8[22] = 8'h6;
    mem8[23] = 8'h7;
    mem8[24] = 8'h8;
    mem8[25] = 8'h9;
    mem8[26] = 8'ha;
    mem8[27] = 8'hb;
    mem8[28] = 8'hc;
    mem8[29] = 8'hd;
    mem8[30] = 8'he;
    mem8[31] = 8'hf;
    mem8[32] = 8'h0;
    mem8[33] = 8'h2;
    mem8[34] = 8'h4;
    mem8[35] = 8'h6;
    mem8[36] = 8'h8;
    mem8[37] = 8'ha;
    mem8[38] = 8'hc;
    mem8[39] = 8'he;
    mem8[40] = 8'h10;
    mem8[41] = 8'h12;
    mem8[42] = 8'h14;
    mem8[43] = 8'h16;
    mem8[44] = 8'h18;
    mem8[45] = 8'h1a;
    mem8[46] = 8'h1c;
    mem8[47] = 8'h1e;
    mem8[48] = 8'h0;
    mem8[49] = 8'h3;
    mem8[50] = 8'h6;
    mem8[51] = 8'h9;
    mem8[52] = 8'hc;
    mem8[53] = 8'hf;
    mem8[54] = 8'h12;
    mem8[55] = 8'h15;
    mem8[56] = 8'h18;
    mem8[57] = 8'h1b;
    mem8[58] = 8'h1e;
    mem8[59] = 8'h21;
    mem8[60] = 8'h24;
    mem8[61] = 8'h27;
    mem8[62] = 8'h2a;
    mem8[63] = 8'h2d;
    mem8[64] = 8'h0;
    mem8[65] = 8'h4;
    mem8[66] = 8'h8;
    mem8[67] = 8'hc;
    mem8[68] = 8'h10;
    mem8[69] = 8'h14;
    mem8[70] = 8'h18;
    mem8[71] = 8'h1c;
    mem8[72] = 8'h20;
    mem8[73] = 8'h24;
    mem8[74] = 8'h28;
    mem8[75] = 8'h2c;
    mem8[76] = 8'h30;
    mem8[77] = 8'h34;
    mem8[78] = 8'h38;
    mem8[79] = 8'h3c;
    mem8[80] = 8'h0;
    mem8[81] = 8'h5;
    mem8[82] = 8'ha;
    mem8[83] = 8'hf;
    mem8[84] = 8'h14;
    mem8[85] = 8'h19;
    mem8[86] = 8'h1e;
    mem8[87] = 8'h23;
    mem8[88] = 8'h28;
    mem8[89] = 8'h2d;
    mem8[90] = 8'h32;
    mem8[91] = 8'h37;
    mem8[92] = 8'h3c;
    mem8[93] = 8'h41;
    mem8[94] = 8'h46;
    mem8[95] = 8'h4b;
    mem8[96] = 8'h0;
    mem8[97] = 8'h6;
    mem8[98] = 8'hc;
    mem8[99] = 8'h12;
    mem8[100] = 8'h18;
    mem8[101] = 8'h1e;
    mem8[102] = 8'h24;
    mem8[103] = 8'h2a;
    mem8[104] = 8'h30;
    mem8[105] = 8'h36;
    mem8[106] = 8'h3c;
    mem8[107] = 8'h42;
    mem8[108] = 8'h48;
    mem8[109] = 8'h4e;
    mem8[110] = 8'h54;
    mem8[111] = 8'h5a;
    mem8[112] = 8'h0;
    mem8[113] = 8'h7;
    mem8[114] = 8'he;
    mem8[115] = 8'h15;
    mem8[116] = 8'h1c;
    mem8[117] = 8'h23;
    mem8[118] = 8'h2a;
    mem8[119] = 8'h31;
    mem8[120] = 8'h38;
    mem8[121] = 8'h3f;
    mem8[122] = 8'h46;
    mem8[123] = 8'h4d;
    mem8[124] = 8'h54;
    mem8[125] = 8'h5b;
    mem8[126] = 8'h62;
    mem8[127] = 8'h69;
    mem8[128] = 8'h0;
    mem8[129] = 8'h8;
    mem8[130] = 8'h10;
    mem8[131] = 8'h18;
    mem8[132] = 8'h20;
    mem8[133] = 8'h28;
    mem8[134] = 8'h30;
    mem8[135] = 8'h38;
    mem8[136] = 8'h40;
    mem8[137] = 8'h48;
    mem8[138] = 8'h50;
    mem8[139] = 8'h58;
    mem8[140] = 8'h60;
    mem8[141] = 8'h68;
    mem8[142] = 8'h70;
    mem8[143] = 8'h78;
    mem8[144] = 8'h0;
    mem8[145] = 8'h9;
    mem8[146] = 8'h12;
    mem8[147] = 8'h1b;
    mem8[148] = 8'h24;
    mem8[149] = 8'h2d;
    mem8[150] = 8'h36;
    mem8[151] = 8'h3f;
    mem8[152] = 8'h48;
    mem8[153] = 8'h51;
    mem8[154] = 8'h5a;
    mem8[155] = 8'h63;
    mem8[156] = 8'h6c;
    mem8[157] = 8'h75;
    mem8[158] = 8'h7e;
    mem8[159] = 8'h87;
    mem8[160] = 8'h0;
    mem8[161] = 8'ha;
    mem8[162] = 8'h14;
    mem8[163] = 8'h1e;
    mem8[164] = 8'h28;
    mem8[165] = 8'h32;
    mem8[166] = 8'h3c;
    mem8[167] = 8'h46;
    mem8[168] = 8'h50;
    mem8[169] = 8'h5a;
    mem8[170] = 8'h64;
    mem8[171] = 8'h6e;
    mem8[172] = 8'h78;
    mem8[173] = 8'h82;
    mem8[174] = 8'h8c;
    mem8[175] = 8'h96;
    mem8[176] = 8'h0;
    mem8[177] = 8'hb;
    mem8[178] = 8'h16;
    mem8[179] = 8'h21;
    mem8[180] = 8'h2c;
    mem8[181] = 8'h37;
    mem8[182] = 8'h42;
    mem8[183] = 8'h4d;
    mem8[184] = 8'h58;
    mem8[185] = 8'h63;
    mem8[186] = 8'h6e;
    mem8[187] = 8'h79;
    mem8[188] = 8'h84;
    mem8[189] = 8'h8f;
    mem8[190] = 8'h9a;
    mem8[191] = 8'ha5;
    mem8[192] = 8'h0;
    mem8[193] = 8'hc;
    mem8[194] = 8'h18;
    mem8[195] = 8'h24;
    mem8[196] = 8'h30;
    mem8[197] = 8'h3c;
    mem8[198] = 8'h48;
    mem8[199] = 8'h54;
    mem8[200] = 8'h60;
    mem8[201] = 8'h6c;
    mem8[202] = 8'h78;
    mem8[203] = 8'h84;
    mem8[204] = 8'h90;
    mem8[205] = 8'h9c;
    mem8[206] = 8'ha8;
    mem8[207] = 8'hb4;
    mem8[208] = 8'h0;
    mem8[209] = 8'hd;
    mem8[210] = 8'h1a;
    mem8[211] = 8'h27;
    mem8[212] = 8'h34;
    mem8[213] = 8'h41;
    mem8[214] = 8'h4e;
    mem8[215] = 8'h5b;
    mem8[216] = 8'h68;
    mem8[217] = 8'h75;
    mem8[218] = 8'h82;
    mem8[219] = 8'h8f;
    mem8[220] = 8'h9c;
    mem8[221] = 8'ha9;
    mem8[222] = 8'hb6;
    mem8[223] = 8'hc3;
    mem8[224] = 8'h0;
    mem8[225] = 8'he;
    mem8[226] = 8'h1c;
    mem8[227] = 8'h2a;
    mem8[228] = 8'h38;
    mem8[229] = 8'h46;
    mem8[230] = 8'h54;
    mem8[231] = 8'h62;
    mem8[232] = 8'h70;
    mem8[233] = 8'h7e;
    mem8[234] = 8'h8c;
    mem8[235] = 8'h9a;
    mem8[236] = 8'ha8;
    mem8[237] = 8'hb6;
    mem8[238] = 8'hc4;
    mem8[239] = 8'hd2;
    mem8[240] = 8'h0;
    mem8[241] = 8'hf;
    mem8[242] = 8'h1e;
    mem8[243] = 8'h2d;
    mem8[244] = 8'h3c;
    mem8[245] = 8'h4b;
    mem8[246] = 8'h5a;
    mem8[247] = 8'h69;
    mem8[248] = 8'h78;
    mem8[249] = 8'h87;
    mem8[250] = 8'h96;
    mem8[251] = 8'ha5;
    mem8[252] = 8'hb4;
    mem8[253] = 8'hc3;
    mem8[254] = 8'hd2;
    mem8[255] = 8'he1;
  end
  assign zext9 = {{4{1'b0}}, io_rhs};
  assign zext11 = {{4{1'b0}}, io_lhs};
  assign sll15 = zext11 << 32'h4;
  assign or17 = sll15 | zext9;

  assign io_out = mem8[or17];

endmodule
