module FastMult(
  input wire[3:0] io_lhs,
  input wire[3:0] io_rhs,
  output wire[7:0] io_out
);
  reg[7:0] mem12[0:255];
  wire[7:0] zext13;
  wire[7:0] zext15;
  wire[7:0] sll19;
  wire[7:0] or21;

  initial begin
    mem12[0] = 8'h0;
    mem12[1] = 8'h0;
    mem12[2] = 8'h0;
    mem12[3] = 8'h0;
    mem12[4] = 8'h0;
    mem12[5] = 8'h0;
    mem12[6] = 8'h0;
    mem12[7] = 8'h0;
    mem12[8] = 8'h0;
    mem12[9] = 8'h0;
    mem12[10] = 8'h0;
    mem12[11] = 8'h0;
    mem12[12] = 8'h0;
    mem12[13] = 8'h0;
    mem12[14] = 8'h0;
    mem12[15] = 8'h0;
    mem12[16] = 8'h0;
    mem12[17] = 8'h1;
    mem12[18] = 8'h2;
    mem12[19] = 8'h3;
    mem12[20] = 8'h4;
    mem12[21] = 8'h5;
    mem12[22] = 8'h6;
    mem12[23] = 8'h7;
    mem12[24] = 8'h8;
    mem12[25] = 8'h9;
    mem12[26] = 8'ha;
    mem12[27] = 8'hb;
    mem12[28] = 8'hc;
    mem12[29] = 8'hd;
    mem12[30] = 8'he;
    mem12[31] = 8'hf;
    mem12[32] = 8'h0;
    mem12[33] = 8'h2;
    mem12[34] = 8'h4;
    mem12[35] = 8'h6;
    mem12[36] = 8'h8;
    mem12[37] = 8'ha;
    mem12[38] = 8'hc;
    mem12[39] = 8'he;
    mem12[40] = 8'h10;
    mem12[41] = 8'h12;
    mem12[42] = 8'h14;
    mem12[43] = 8'h16;
    mem12[44] = 8'h18;
    mem12[45] = 8'h1a;
    mem12[46] = 8'h1c;
    mem12[47] = 8'h1e;
    mem12[48] = 8'h0;
    mem12[49] = 8'h3;
    mem12[50] = 8'h6;
    mem12[51] = 8'h9;
    mem12[52] = 8'hc;
    mem12[53] = 8'hf;
    mem12[54] = 8'h12;
    mem12[55] = 8'h15;
    mem12[56] = 8'h18;
    mem12[57] = 8'h1b;
    mem12[58] = 8'h1e;
    mem12[59] = 8'h21;
    mem12[60] = 8'h24;
    mem12[61] = 8'h27;
    mem12[62] = 8'h2a;
    mem12[63] = 8'h2d;
    mem12[64] = 8'h0;
    mem12[65] = 8'h4;
    mem12[66] = 8'h8;
    mem12[67] = 8'hc;
    mem12[68] = 8'h10;
    mem12[69] = 8'h14;
    mem12[70] = 8'h18;
    mem12[71] = 8'h1c;
    mem12[72] = 8'h20;
    mem12[73] = 8'h24;
    mem12[74] = 8'h28;
    mem12[75] = 8'h2c;
    mem12[76] = 8'h30;
    mem12[77] = 8'h34;
    mem12[78] = 8'h38;
    mem12[79] = 8'h3c;
    mem12[80] = 8'h0;
    mem12[81] = 8'h5;
    mem12[82] = 8'ha;
    mem12[83] = 8'hf;
    mem12[84] = 8'h14;
    mem12[85] = 8'h19;
    mem12[86] = 8'h1e;
    mem12[87] = 8'h23;
    mem12[88] = 8'h28;
    mem12[89] = 8'h2d;
    mem12[90] = 8'h32;
    mem12[91] = 8'h37;
    mem12[92] = 8'h3c;
    mem12[93] = 8'h41;
    mem12[94] = 8'h46;
    mem12[95] = 8'h4b;
    mem12[96] = 8'h0;
    mem12[97] = 8'h6;
    mem12[98] = 8'hc;
    mem12[99] = 8'h12;
    mem12[100] = 8'h18;
    mem12[101] = 8'h1e;
    mem12[102] = 8'h24;
    mem12[103] = 8'h2a;
    mem12[104] = 8'h30;
    mem12[105] = 8'h36;
    mem12[106] = 8'h3c;
    mem12[107] = 8'h42;
    mem12[108] = 8'h48;
    mem12[109] = 8'h4e;
    mem12[110] = 8'h54;
    mem12[111] = 8'h5a;
    mem12[112] = 8'h0;
    mem12[113] = 8'h7;
    mem12[114] = 8'he;
    mem12[115] = 8'h15;
    mem12[116] = 8'h1c;
    mem12[117] = 8'h23;
    mem12[118] = 8'h2a;
    mem12[119] = 8'h31;
    mem12[120] = 8'h38;
    mem12[121] = 8'h3f;
    mem12[122] = 8'h46;
    mem12[123] = 8'h4d;
    mem12[124] = 8'h54;
    mem12[125] = 8'h5b;
    mem12[126] = 8'h62;
    mem12[127] = 8'h69;
    mem12[128] = 8'h0;
    mem12[129] = 8'h8;
    mem12[130] = 8'h10;
    mem12[131] = 8'h18;
    mem12[132] = 8'h20;
    mem12[133] = 8'h28;
    mem12[134] = 8'h30;
    mem12[135] = 8'h38;
    mem12[136] = 8'h40;
    mem12[137] = 8'h48;
    mem12[138] = 8'h50;
    mem12[139] = 8'h58;
    mem12[140] = 8'h60;
    mem12[141] = 8'h68;
    mem12[142] = 8'h70;
    mem12[143] = 8'h78;
    mem12[144] = 8'h0;
    mem12[145] = 8'h9;
    mem12[146] = 8'h12;
    mem12[147] = 8'h1b;
    mem12[148] = 8'h24;
    mem12[149] = 8'h2d;
    mem12[150] = 8'h36;
    mem12[151] = 8'h3f;
    mem12[152] = 8'h48;
    mem12[153] = 8'h51;
    mem12[154] = 8'h5a;
    mem12[155] = 8'h63;
    mem12[156] = 8'h6c;
    mem12[157] = 8'h75;
    mem12[158] = 8'h7e;
    mem12[159] = 8'h87;
    mem12[160] = 8'h0;
    mem12[161] = 8'ha;
    mem12[162] = 8'h14;
    mem12[163] = 8'h1e;
    mem12[164] = 8'h28;
    mem12[165] = 8'h32;
    mem12[166] = 8'h3c;
    mem12[167] = 8'h46;
    mem12[168] = 8'h50;
    mem12[169] = 8'h5a;
    mem12[170] = 8'h64;
    mem12[171] = 8'h6e;
    mem12[172] = 8'h78;
    mem12[173] = 8'h82;
    mem12[174] = 8'h8c;
    mem12[175] = 8'h96;
    mem12[176] = 8'h0;
    mem12[177] = 8'hb;
    mem12[178] = 8'h16;
    mem12[179] = 8'h21;
    mem12[180] = 8'h2c;
    mem12[181] = 8'h37;
    mem12[182] = 8'h42;
    mem12[183] = 8'h4d;
    mem12[184] = 8'h58;
    mem12[185] = 8'h63;
    mem12[186] = 8'h6e;
    mem12[187] = 8'h79;
    mem12[188] = 8'h84;
    mem12[189] = 8'h8f;
    mem12[190] = 8'h9a;
    mem12[191] = 8'ha5;
    mem12[192] = 8'h0;
    mem12[193] = 8'hc;
    mem12[194] = 8'h18;
    mem12[195] = 8'h24;
    mem12[196] = 8'h30;
    mem12[197] = 8'h3c;
    mem12[198] = 8'h48;
    mem12[199] = 8'h54;
    mem12[200] = 8'h60;
    mem12[201] = 8'h6c;
    mem12[202] = 8'h78;
    mem12[203] = 8'h84;
    mem12[204] = 8'h90;
    mem12[205] = 8'h9c;
    mem12[206] = 8'ha8;
    mem12[207] = 8'hb4;
    mem12[208] = 8'h0;
    mem12[209] = 8'hd;
    mem12[210] = 8'h1a;
    mem12[211] = 8'h27;
    mem12[212] = 8'h34;
    mem12[213] = 8'h41;
    mem12[214] = 8'h4e;
    mem12[215] = 8'h5b;
    mem12[216] = 8'h68;
    mem12[217] = 8'h75;
    mem12[218] = 8'h82;
    mem12[219] = 8'h8f;
    mem12[220] = 8'h9c;
    mem12[221] = 8'ha9;
    mem12[222] = 8'hb6;
    mem12[223] = 8'hc3;
    mem12[224] = 8'h0;
    mem12[225] = 8'he;
    mem12[226] = 8'h1c;
    mem12[227] = 8'h2a;
    mem12[228] = 8'h38;
    mem12[229] = 8'h46;
    mem12[230] = 8'h54;
    mem12[231] = 8'h62;
    mem12[232] = 8'h70;
    mem12[233] = 8'h7e;
    mem12[234] = 8'h8c;
    mem12[235] = 8'h9a;
    mem12[236] = 8'ha8;
    mem12[237] = 8'hb6;
    mem12[238] = 8'hc4;
    mem12[239] = 8'hd2;
    mem12[240] = 8'h0;
    mem12[241] = 8'hf;
    mem12[242] = 8'h1e;
    mem12[243] = 8'h2d;
    mem12[244] = 8'h3c;
    mem12[245] = 8'h4b;
    mem12[246] = 8'h5a;
    mem12[247] = 8'h69;
    mem12[248] = 8'h78;
    mem12[249] = 8'h87;
    mem12[250] = 8'h96;
    mem12[251] = 8'ha5;
    mem12[252] = 8'hb4;
    mem12[253] = 8'hc3;
    mem12[254] = 8'hd2;
    mem12[255] = 8'he1;
  end
  assign zext13 = {{4{1'b0}}, io_rhs};
  assign zext15 = {{4{1'b0}}, io_lhs};
  assign sll19 = zext15 << 32'h4;
  assign or21 = sll19 | zext13;

  assign io_out = mem12[or21];

endmodule
