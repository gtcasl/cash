module FastMult(
  input wire[3:0] io_lhs,
  input wire[3:0] io_rhs,
  output wire[7:0] io_out
);
  wire[7:0] zext17;
  wire[7:0] zext15;
  wire[7:0] sll21;
  wire[7:0] or23;
  reg[7:0] mem14[0:255];

  assign zext17 = {{4{1'b0}}, io_lhs};
  assign zext15 = {{4{1'b0}}, io_rhs};
  assign sll21 = zext17 << 32'h4;
  assign or23 = sll21 | zext15;
  initial begin
    mem14[0] = 8'h0;
    mem14[1] = 8'h0;
    mem14[2] = 8'h0;
    mem14[3] = 8'h0;
    mem14[4] = 8'h0;
    mem14[5] = 8'h0;
    mem14[6] = 8'h0;
    mem14[7] = 8'h0;
    mem14[8] = 8'h0;
    mem14[9] = 8'h0;
    mem14[10] = 8'h0;
    mem14[11] = 8'h0;
    mem14[12] = 8'h0;
    mem14[13] = 8'h0;
    mem14[14] = 8'h0;
    mem14[15] = 8'h0;
    mem14[16] = 8'h0;
    mem14[17] = 8'h1;
    mem14[18] = 8'h2;
    mem14[19] = 8'h3;
    mem14[20] = 8'h4;
    mem14[21] = 8'h5;
    mem14[22] = 8'h6;
    mem14[23] = 8'h7;
    mem14[24] = 8'h8;
    mem14[25] = 8'h9;
    mem14[26] = 8'ha;
    mem14[27] = 8'hb;
    mem14[28] = 8'hc;
    mem14[29] = 8'hd;
    mem14[30] = 8'he;
    mem14[31] = 8'hf;
    mem14[32] = 8'h0;
    mem14[33] = 8'h2;
    mem14[34] = 8'h4;
    mem14[35] = 8'h6;
    mem14[36] = 8'h8;
    mem14[37] = 8'ha;
    mem14[38] = 8'hc;
    mem14[39] = 8'he;
    mem14[40] = 8'h10;
    mem14[41] = 8'h12;
    mem14[42] = 8'h14;
    mem14[43] = 8'h16;
    mem14[44] = 8'h18;
    mem14[45] = 8'h1a;
    mem14[46] = 8'h1c;
    mem14[47] = 8'h1e;
    mem14[48] = 8'h0;
    mem14[49] = 8'h3;
    mem14[50] = 8'h6;
    mem14[51] = 8'h9;
    mem14[52] = 8'hc;
    mem14[53] = 8'hf;
    mem14[54] = 8'h12;
    mem14[55] = 8'h15;
    mem14[56] = 8'h18;
    mem14[57] = 8'h1b;
    mem14[58] = 8'h1e;
    mem14[59] = 8'h21;
    mem14[60] = 8'h24;
    mem14[61] = 8'h27;
    mem14[62] = 8'h2a;
    mem14[63] = 8'h2d;
    mem14[64] = 8'h0;
    mem14[65] = 8'h4;
    mem14[66] = 8'h8;
    mem14[67] = 8'hc;
    mem14[68] = 8'h10;
    mem14[69] = 8'h14;
    mem14[70] = 8'h18;
    mem14[71] = 8'h1c;
    mem14[72] = 8'h20;
    mem14[73] = 8'h24;
    mem14[74] = 8'h28;
    mem14[75] = 8'h2c;
    mem14[76] = 8'h30;
    mem14[77] = 8'h34;
    mem14[78] = 8'h38;
    mem14[79] = 8'h3c;
    mem14[80] = 8'h0;
    mem14[81] = 8'h5;
    mem14[82] = 8'ha;
    mem14[83] = 8'hf;
    mem14[84] = 8'h14;
    mem14[85] = 8'h19;
    mem14[86] = 8'h1e;
    mem14[87] = 8'h23;
    mem14[88] = 8'h28;
    mem14[89] = 8'h2d;
    mem14[90] = 8'h32;
    mem14[91] = 8'h37;
    mem14[92] = 8'h3c;
    mem14[93] = 8'h41;
    mem14[94] = 8'h46;
    mem14[95] = 8'h4b;
    mem14[96] = 8'h0;
    mem14[97] = 8'h6;
    mem14[98] = 8'hc;
    mem14[99] = 8'h12;
    mem14[100] = 8'h18;
    mem14[101] = 8'h1e;
    mem14[102] = 8'h24;
    mem14[103] = 8'h2a;
    mem14[104] = 8'h30;
    mem14[105] = 8'h36;
    mem14[106] = 8'h3c;
    mem14[107] = 8'h42;
    mem14[108] = 8'h48;
    mem14[109] = 8'h4e;
    mem14[110] = 8'h54;
    mem14[111] = 8'h5a;
    mem14[112] = 8'h0;
    mem14[113] = 8'h7;
    mem14[114] = 8'he;
    mem14[115] = 8'h15;
    mem14[116] = 8'h1c;
    mem14[117] = 8'h23;
    mem14[118] = 8'h2a;
    mem14[119] = 8'h31;
    mem14[120] = 8'h38;
    mem14[121] = 8'h3f;
    mem14[122] = 8'h46;
    mem14[123] = 8'h4d;
    mem14[124] = 8'h54;
    mem14[125] = 8'h5b;
    mem14[126] = 8'h62;
    mem14[127] = 8'h69;
    mem14[128] = 8'h0;
    mem14[129] = 8'h8;
    mem14[130] = 8'h10;
    mem14[131] = 8'h18;
    mem14[132] = 8'h20;
    mem14[133] = 8'h28;
    mem14[134] = 8'h30;
    mem14[135] = 8'h38;
    mem14[136] = 8'h40;
    mem14[137] = 8'h48;
    mem14[138] = 8'h50;
    mem14[139] = 8'h58;
    mem14[140] = 8'h60;
    mem14[141] = 8'h68;
    mem14[142] = 8'h70;
    mem14[143] = 8'h78;
    mem14[144] = 8'h0;
    mem14[145] = 8'h9;
    mem14[146] = 8'h12;
    mem14[147] = 8'h1b;
    mem14[148] = 8'h24;
    mem14[149] = 8'h2d;
    mem14[150] = 8'h36;
    mem14[151] = 8'h3f;
    mem14[152] = 8'h48;
    mem14[153] = 8'h51;
    mem14[154] = 8'h5a;
    mem14[155] = 8'h63;
    mem14[156] = 8'h6c;
    mem14[157] = 8'h75;
    mem14[158] = 8'h7e;
    mem14[159] = 8'h87;
    mem14[160] = 8'h0;
    mem14[161] = 8'ha;
    mem14[162] = 8'h14;
    mem14[163] = 8'h1e;
    mem14[164] = 8'h28;
    mem14[165] = 8'h32;
    mem14[166] = 8'h3c;
    mem14[167] = 8'h46;
    mem14[168] = 8'h50;
    mem14[169] = 8'h5a;
    mem14[170] = 8'h64;
    mem14[171] = 8'h6e;
    mem14[172] = 8'h78;
    mem14[173] = 8'h82;
    mem14[174] = 8'h8c;
    mem14[175] = 8'h96;
    mem14[176] = 8'h0;
    mem14[177] = 8'hb;
    mem14[178] = 8'h16;
    mem14[179] = 8'h21;
    mem14[180] = 8'h2c;
    mem14[181] = 8'h37;
    mem14[182] = 8'h42;
    mem14[183] = 8'h4d;
    mem14[184] = 8'h58;
    mem14[185] = 8'h63;
    mem14[186] = 8'h6e;
    mem14[187] = 8'h79;
    mem14[188] = 8'h84;
    mem14[189] = 8'h8f;
    mem14[190] = 8'h9a;
    mem14[191] = 8'ha5;
    mem14[192] = 8'h0;
    mem14[193] = 8'hc;
    mem14[194] = 8'h18;
    mem14[195] = 8'h24;
    mem14[196] = 8'h30;
    mem14[197] = 8'h3c;
    mem14[198] = 8'h48;
    mem14[199] = 8'h54;
    mem14[200] = 8'h60;
    mem14[201] = 8'h6c;
    mem14[202] = 8'h78;
    mem14[203] = 8'h84;
    mem14[204] = 8'h90;
    mem14[205] = 8'h9c;
    mem14[206] = 8'ha8;
    mem14[207] = 8'hb4;
    mem14[208] = 8'h0;
    mem14[209] = 8'hd;
    mem14[210] = 8'h1a;
    mem14[211] = 8'h27;
    mem14[212] = 8'h34;
    mem14[213] = 8'h41;
    mem14[214] = 8'h4e;
    mem14[215] = 8'h5b;
    mem14[216] = 8'h68;
    mem14[217] = 8'h75;
    mem14[218] = 8'h82;
    mem14[219] = 8'h8f;
    mem14[220] = 8'h9c;
    mem14[221] = 8'ha9;
    mem14[222] = 8'hb6;
    mem14[223] = 8'hc3;
    mem14[224] = 8'h0;
    mem14[225] = 8'he;
    mem14[226] = 8'h1c;
    mem14[227] = 8'h2a;
    mem14[228] = 8'h38;
    mem14[229] = 8'h46;
    mem14[230] = 8'h54;
    mem14[231] = 8'h62;
    mem14[232] = 8'h70;
    mem14[233] = 8'h7e;
    mem14[234] = 8'h8c;
    mem14[235] = 8'h9a;
    mem14[236] = 8'ha8;
    mem14[237] = 8'hb6;
    mem14[238] = 8'hc4;
    mem14[239] = 8'hd2;
    mem14[240] = 8'h0;
    mem14[241] = 8'hf;
    mem14[242] = 8'h1e;
    mem14[243] = 8'h2d;
    mem14[244] = 8'h3c;
    mem14[245] = 8'h4b;
    mem14[246] = 8'h5a;
    mem14[247] = 8'h69;
    mem14[248] = 8'h78;
    mem14[249] = 8'h87;
    mem14[250] = 8'h96;
    mem14[251] = 8'ha5;
    mem14[252] = 8'hb4;
    mem14[253] = 8'hc3;
    mem14[254] = 8'hd2;
    mem14[255] = 8'he1;
  end

  assign io_out = mem14[or23];

endmodule
